// =============================================================
// Definitions for Virtual USB code in Modelsim
//
// Copyright (c) 2023 Simon Southwell.
//
// This file is part of usbModel pattern generator.
//
// This code is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
//
// The code is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this code. If not, see <http://www.gnu.org/licenses/>.
//
// =============================================================

`ifndef _USB_VH_
`define _USB_VH_

`define NODE_NUM               0
`define CLKCOUNT               1
`define RESET_STATE            2
`define PULLUP                 3
`define OUTEN                  4
`define LINE                   5

`define UVH_STOP               1001
`define UVH_FINISH             1002

`endif